module top_module (vec,outv, o2,o1,o0 );
input [2:0] vec;
output o2,o1,o0;
output [2:0] outv;

assign outv= vec;
assign o2= vec[2]; 
assign o1= vec[1]; 
assign o0= vec[0]; 

endmodule
