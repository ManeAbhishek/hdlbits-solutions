module top_module(
    input a,
    input b,
    input c,
    input d,
    output out,
    output out_n ); 
wire x; wire y ; wire z;
    and(x,a,b);
    and(y,c,d);
    or(z,x,y);
    assign out = z;
    assign out_n = ~z;
    


endmodule
